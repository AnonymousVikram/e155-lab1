../src/lab1_vk.sv